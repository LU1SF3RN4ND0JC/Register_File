library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity decoder5x32 is
    Port ( inp : in  STD_LOGIC_VECTOR (4 downto 0);
           outp : out  STD_LOGIC_VECTOR (31 downto 0));
end decoder5x32;

architecture decoder_arch of decoder5x32 is

begin
outp <= "00000000000000000000000000000001" when inp = "00000" else
		"00000000000000000000000000000010" when inp = "00001" else
		"00000000000000000000000000000100" when inp = "00010" else
		"00000000000000000000000000001000" when inp = "00011" else
		"00000000000000000000000000010000" when inp = "00100" else
		"00000000000000000000000000100000" when inp = "00101" else
		"00000000000000000000000001000000" when inp = "00110" else
		"00000000000000000000000010000000" when inp = "00111" else
		"00000000000000000000000100000000" when inp = "01000" else
		"00000000000000000000001000000000" when inp = "01001" else
		"00000000000000000000010000000000" when inp = "01010" else
		"00000000000000000000100000000000" when inp = "01011" else
		"00000000000000000001000000000000" when inp = "01100" else
		"00000000000000000010000000000000" when inp = "01101" else
		"00000000000000000100000000000000" when inp = "01110" else
		"00000000000000001000000000000000" when inp = "01111" else
		"00000000000000010000000000000000" when inp = "10000" else
		"00000000000000100000000000000000" when inp = "10001" else
		"00000000000001000000000000000000" when inp = "10010" else
		"00000000000010000000000000000000" when inp = "10011" else
		"00000000000100000000000000000000" when inp = "10100" else
		"00000000001000000000000000000000" when inp = "10101" else
		"00000000010000000000000000000000" when inp = "10110" else
		"00000000100000000000000000000000" when inp = "10111" else
		"00000001000000000000000000000000" when inp = "11000" else
		"00000010000000000000000000000000" when inp = "11001" else
		"00000100000000000000000000000000" when inp = "11010" else
		"00001000000000000000000000000000" when inp = "11011" else
		"00010000000000000000000000000000" when inp = "11100" else
		"00100000000000000000000000000000" when inp = "11101" else
		"01000000000000000000000000000000" when inp = "11110" else
		"10000000000000000000000000000000" when inp = "11111" else
		"ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ" ;
end decoder_arch;