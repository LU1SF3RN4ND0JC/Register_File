library ieee;
use ieee.std_logic_1164.all;

entity mux5x32_tb is 
end mux5x32_tb;

architecture mux_tb of mux5x32_tb is
    component mux5x32
        port(
            I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,I16,I17,I18,I19,I20,I21,I22,I23,I24,I25,I26,I27,I28,I29,I30,I31 : in  STD_LOGIC_VECTOR (31 downto 0);
            Selector : in  STD_LOGIC_VECTOR (4 downto 0);
            O : out  STD_LOGIC_VECTOR (31 downto 0)
        );
    end component;
        signal t_I0,t_I1,t_I2,t_I3,t_I4,t_I5,t_I6,t_I7,t_I8,t_I9,t_I10,t_I11,t_I12,t_I13,t_I14,t_I15,t_I16,t_I17,t_I18,t_I19,t_I20,t_I21,t_I22,t_I23,t_I24,t_I25,t_I26,t_I27,t_I28,t_I29,t_I30,t_I31 : STD_LOGIC_VECTOR (31 downto 0);
        signal t_Selector : STD_LOGIC_VECTOR (4 downto 0);
        signal t_O : STD_LOGIC_VECTOR (31 downto 0);
    begin
        uut: mux5x32 port map(Selector=>t_Selector,O=>t_O,I0=>t_I0,I1=>t_I1,I2=>t_I2,I3=>t_I3,I4=>t_I4,I5=>t_I5,I6=>t_I6,I7=>t_I7,I8=>t_I8,I9=>t_I9,I10=>t_I10,I11=>t_I11,I12=>t_I12,I13=>t_I13,I14=>t_I14,I15=>t_I15,I16=>t_I16,I17=>t_I17,I18=>t_I18,I19=>t_I19,I20=>t_I20,I21=>t_I21,I22=>t_I22,I23=>t_I23,I24=>t_I24,I25=>t_I25,I26=>t_I26,I27=>t_I27,I28=>t_I28,I29=>t_I29,I30=>t_I30,I31=>t_I31);

    process
    begin 
        t_I0<= "11111111111111111111111111111111";
        t_I1<= "11111111111111111111111111111110";
        t_I2<= "11111111111111111111111111111111";
        t_I3<= "11111111111111111111111111111110";
        t_I4<= "11111111111111111111111111111111";
        t_I5<= "11111111111111111111111111111110";
        t_I6<= "11111111111111111111111111111111";
        t_I7<= "11111111111111111111111111111111";
        t_I8<= "11111111111111111111111111111110";
        t_I9<= "11111111111111111111111111111111";
        t_I10<= "11111111111111111111111111111110";
        t_I11<= "11111111111111111111111111111111";
        t_I12<= "11111111111111111111111111111110";
        t_I13<= "11111111111111111111111111111111";
        t_I14<= "11111111111111111111111111111111";
        t_I15<= "11111111111111111111111111111111";
        t_I16<= "11111111111111111111111111111111";
        t_I17<= "11111111111111111111111111111111";
        t_I18<= "11111111111111111111111111111111";
        t_I19<= "11111111111111111111111111111111";
        t_I20<= "11111111111111111111111111111111";
        t_I21<= "11111111111111111111111111111111";
        t_I22<= "11111111111111111111111111111111";
        t_I23<= "11111111111111111111111111111111";
        t_I24<= "11111111111111111111111111111111";
        t_I25<= "11111111111111111111111111111111";
        t_I26<= "11111111111111111111111111111111";
        t_I27<= "11111111111111111111111111111111";
        t_I28<= "11111111111111111111111111111111";
        t_I29<= "11111111111111111111111111111111";
        t_I30<= "11111111111111111111111111111111";
        t_I31<= "00000000000000000000000000000000"; 
        t_selector <= "11111";
        wait for 200 ns;
        t_I0<= "00111111111111111111111111111100";
        t_I1<= "11111111111111111111111111111110";
        t_I2<= "11111111111111111111111111111111";
        t_I3<= "11111111111111111111111111111110";
        t_I4<= "11111111111111111111111111111111";
        t_I5<= "11111111111111111111111111111110";
        t_I6<= "11111111111111111111111111111111";
        t_I7<= "11111111111111111111111111111111";
        t_I8<= "11111111111111111111111111111110";
        t_I9<= "11111111111111111111111111111111";
        t_I10<= "11111111111111111111111111111110";
        t_I11<= "11111111111111111111111111111111";
        t_I12<= "11111111111111111111111111111110";
        t_I13<= "11111111111111111111111111111111";
        t_I14<= "11111111111111111111111111111111";
        t_I15<= "11111111111111111111111111111111";
        t_I16<= "11111111111111111111111111111111";
        t_I17<= "11111111111111111111111111111111";
        t_I18<= "11111111111111111111111111111111";
        t_I19<= "11111111111111111111111111111111";
        t_I20<= "11111111111111111111111111111111";
        t_I21<= "11111111111111111111111111111111";
        t_I22<= "11111111111111111111111111111111";
        t_I23<= "11111111111111111111111111111111";
        t_I24<= "11111111111111111111111111111111";
        t_I25<= "11111111111111111111111111111111";
        t_I26<= "11111111111111111111111111111111";
        t_I27<= "11111111111111111111111111111111";
        t_I28<= "11111111111111111111111111111111";
        t_I29<= "11111111111111111111111111111111";
        t_I30<= "11111111111111111111111111111111";
        t_I31<= "00000000000000000000000000000000";
        t_selector <= "00000";
        wait for 200 ns;
    end process;

end mux_tb;